abcDEF
\a@3jja_=\ 
