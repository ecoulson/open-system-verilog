          




