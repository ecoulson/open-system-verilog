          



        
