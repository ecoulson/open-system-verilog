"foo"
"bar\""
"bar\n"
"fail!
