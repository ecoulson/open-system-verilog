+ - ! ~ & ~& | ~| ^ ~^ ^~ ++ -- ** * / %
>> << >>> <<< < <= > >= inside dist == != === !==
==? !=? && || -> <-> = += -= *= /= %= &= ^= |=
<<= >>= <<<= >>>=
