// A comment
// Another one
/*
*
* BLOCK
* COMMENT
*
*/
