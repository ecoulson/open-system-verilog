"foo"
"bar\""
"bar\n"
"A
Long
Long
Long
Boi"
"fail!
