@#$()[]{};:',.?`_\
